import ALU::*;

(* synthesize *)
module mkALUTests(Empty);
    rule test;
        $display("mkALUTests running...");
        $finish();
    endrule
endmodule
