typedef Bit#(32) Word;
typedef Word ProgramCounter;
typedef Bit#(5) RegisterIndex;
